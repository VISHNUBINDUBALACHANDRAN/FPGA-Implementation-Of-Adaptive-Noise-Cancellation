Library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use IEEE.numeric_std.all;
USE STD.TEXTIO.ALL;

Entity FIR_TB is 
  generic ( n : integer := 16;nn : integer := 32; tab:integer:=50; samples:integer:=5000);
  port(   clk:in std_logic;
        FIRin:inout std_logic_vector(n-1 downto 0):=(others=>'0');
        FIRout:inout std_logic_vector((2*n)-1 downto 0);
        FIRout1:inout std_logic_vector((2*n)-1 downto 0));
end entity;

Architecture test_bench of FIR_TB is 

component FIR_filter is
  generic ( n : integer := 16; tab:integer:=50);
    port(clk:in  std_logic;
           x:in  std_logic_vector(n-1 downto 0);
           y:out std_logic_vector((2*n)-1 downto 0)
         );
end component;

component FIR_filterm_32 is
  generic ( n : integer := 32; tab:integer:=50);
    port(clk:in  std_logic;
           x:in  std_logic_vector(n-1 downto 0);
           y:out std_logic_vector((2*n)-1 downto 0)
         );
end component;


type signalType is array (1 to samples) of std_logic_vector(n-1 downto 0);
type signalType1 is array (1 to samples) of std_logic_vector(31 downto 0);

type signalTypeInt is array (1 to samples) of integer;
signal input:signalType;
signal input1:signalType1;
signal count:integer:=1;
signal ss,ss1:integer:=0;
signal FIRde,fir_er: std_logic_vector(31 downto 0):=(others=>'0');
signal ps: std_logic_vector(15 downto 0):=(others=>'0');
signal ec:integer:=65536;
  begin
   process(clk)
     
     variable sig,sig1:signalTypeInt;
     variable pp:integer;
     
    file text_var:text;
    variable line_var:line;
    variable std_logic_vec:std_logic_vector(7 downto 0);
     begin
   if rising_edge(clk) then 
        file_open(text_var,"ECG_IN.txt",read_mode);
        for i in 1 to samples loop
           if(NOT ENDFILE(text_var))then
              readline(text_var,line_var);
              read(line_var,sig(i));       
             input(i)<=std_logic_vector(to_signed(sig(i),n)); 
             end if;
          end loop;
        file_close(text_var);
        
        
        file_open(text_var,"ECG_de.txt",read_mode);
        for i in 1 to samples loop
           if(NOT ENDFILE(text_var))then
              readline(text_var,line_var);
              read(line_var,sig1(i));   
              pp:=(sig1(i) * 10000) ;   
             input1(i)<=std_logic_vector(to_signed(pp,32)); 
             end if;
          end loop;
        file_close(text_var);
        
        
          
          count<=count+1;
           if count>=samples then
             count<=1;
           end if;  
     end if;
   end process;
  
  FIRin<=input(count);
  
  FIR:FIR_filter generic map(n,tab)
            port map(clk,FIRin,FIRout);
            
  FIRde<=input1(count);
  
fir_er<= (FIRout - FIRde);

ss<= ((conv_integer(fir_er))/ec);

ps<= std_logic_vector(to_signed(ss,16));

  FIR1:FIR_filter generic map(n,tab)
            port map(clk,ps,FIRout1);



end;
  